-------------------------------------------------------------------------------
--                                                                           --
-- CERN BE-CO-HT         GN4124 core for PCIe FMC carrier                    --
--                       http://www.ohwr.org/projects/gn4124-core            --
-------------------------------------------------------------------------------
--
-- unit name: GN4124 core arbiter (arbiter.vhd)
--
-- authors: Simon Deprez (simon.deprez@cern.ch)
--          Matthieu Cattin (matthieu.cattin@cern.ch)
--
-- date: 12-08-2010
--
-- version: 0.1
--
-- description: Arbitrates PCIe accesses between Wishbone master,
--              L2P DMA master and P2L DMA master
--
-- dependencies:
--
-------------------------------------------------------------------------------
-- last changes: 23-09-2010 (mcattin) Add FF on data path and
--                                    change valid request logic
-------------------------------------------------------------------------------
-- TODO: -
--       -
--       -
-------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
use work.gn4124_core_pkg.all;


entity arbiter is
  port
    (
      ---------------------------------------------------------
      -- Clock/Reset
      clk_i   : in std_logic;
      rst_n_i : in std_logic;

      ---------------------------------------------------------
      -- From Wishbone master (wbm) to arbiter (arb)
      wbm_arb_valid_i  : in  std_logic;
      wbm_arb_dframe_i : in  std_logic;
      wbm_arb_data_i   : in  std_logic_vector(31 downto 0);
      wbm_arb_req_i    : in  std_logic;
      arb_wbm_gnt_o    : out std_logic;

      ---------------------------------------------------------
      -- From DMA pdmuencer (pdm) to arbiter (arb)
      pdm_arb_valid_i  : in  std_logic;
      pdm_arb_dframe_i : in  std_logic;
      pdm_arb_data_i   : in  std_logic_vector(31 downto 0);
      pdm_arb_req_i    : in  std_logic;
      arb_pdm_gnt_o    : out std_logic;

      ---------------------------------------------------------
      -- From P2L DMA master (ldm) to arbiter (arb)
      ldm_arb_valid_i  : in  std_logic;
      ldm_arb_dframe_i : in  std_logic;
      ldm_arb_data_i   : in  std_logic_vector(31 downto 0);
      ldm_arb_req_i    : in  std_logic;
      arb_ldm_gnt_o    : out std_logic;

      ---------------------------------------------------------
      -- From arbiter (arb) to serializer (ser)
      arb_ser_valid_o  : out std_logic;
      arb_ser_dframe_o : out std_logic;
      arb_ser_data_o   : out std_logic_vector(31 downto 0)
      );
end arbiter;


architecture behaviour of arbiter is


---------------------------------------------------------
  -- Signal declarations
  signal wbm_arb_req_valid : std_logic;
  signal pdm_arb_req_valid : std_logic;
  signal ldm_arb_req_valid : std_logic;
  signal arb_wbm_gnt       : std_logic;
  signal arb_pdm_gnt       : std_logic;
  signal arb_ldm_gnt       : std_logic;
  signal eop               : std_logic;  -- End of packet


begin


  -- A request is valid only if the access not already granted to another source
  wbm_arb_req_valid <= wbm_arb_req_i and (not(arb_pdm_gnt) and not(arb_ldm_gnt));
  pdm_arb_req_valid <= pdm_arb_req_i and (not(arb_wbm_gnt) and not(arb_ldm_gnt));
  ldm_arb_req_valid <= ldm_arb_req_i and (not(arb_wbm_gnt) and not(arb_pdm_gnt));

  -- Detect end of packet to delimit the arbitration phase
  eop <= ((arb_wbm_gnt and not(wbm_arb_dframe_i) and wbm_arb_valid_i) or
          (arb_pdm_gnt and not(pdm_arb_dframe_i) and pdm_arb_valid_i) or
          (arb_ldm_gnt and not(ldm_arb_dframe_i) and ldm_arb_valid_i));

  -----------------------------------------------------------------------------
  -- Arbitration is started when a valid request is present and ends when the
  -- EOP condition is detected
  --
  -- Strict priority arbitration scheme
  -- Highest : WBM request
  --         : LDM request
  -- Lowest  : PDM request
  -----------------------------------------------------------------------------
  process (clk_i, rst_n_i)
  begin
    if(rst_n_i = c_RST_ACTIVE) then
      arb_wbm_gnt <= '0';
      arb_pdm_gnt <= '0';
      arb_ldm_gnt <= '0';
    elsif rising_edge(clk_i) then
      --if (arb_req_valid = '1') then
      if (wbm_arb_req_valid = '1') then
        arb_wbm_gnt <= '1';
        arb_pdm_gnt <= '0';
        arb_ldm_gnt <= '0';
      elsif (ldm_arb_req_valid = '1') then
        arb_wbm_gnt <= '0';
        arb_pdm_gnt <= '0';
        arb_ldm_gnt <= '1';
      elsif (pdm_arb_req_valid = '1') then
        arb_wbm_gnt <= '0';
        arb_pdm_gnt <= '1';
        arb_ldm_gnt <= '0';
      elsif (eop = '1') then
        arb_wbm_gnt <= '0';
        arb_pdm_gnt <= '0';
        arb_ldm_gnt <= '0';
      end if;
    end if;
  end process;

  process (clk_i, rst_n_i)
  begin
    if rst_n_i = '0' then
      arb_ser_valid_o  <= '0';
      arb_ser_dframe_o <= '0';
      arb_ser_data_o   <= (others => '0');
    elsif rising_edge(clk_i) then
      if arb_wbm_gnt = '1' then
        arb_ser_valid_o  <= wbm_arb_valid_i;
        arb_ser_dframe_o <= wbm_arb_dframe_i;
        arb_ser_data_o   <= wbm_arb_data_i;
      elsif arb_pdm_gnt = '1' then
        arb_ser_valid_o  <= pdm_arb_valid_i;
        arb_ser_dframe_o <= pdm_arb_dframe_i;
        arb_ser_data_o   <= pdm_arb_data_i;
      elsif arb_ldm_gnt = '1' then
        arb_ser_valid_o  <= ldm_arb_valid_i;
        arb_ser_dframe_o <= ldm_arb_dframe_i;
        arb_ser_data_o   <= ldm_arb_data_i;
      else
        arb_ser_valid_o  <= '0';
        arb_ser_dframe_o <= '0';
        arb_ser_data_o   <= (others => '0');
      end if;
    end if;
  end process;

  arb_wbm_gnt_o <= arb_wbm_gnt;
  arb_pdm_gnt_o <= arb_pdm_gnt;
  arb_ldm_gnt_o <= arb_ldm_gnt;

end behaviour;
