--------------------------------------------------------------------------------
--                                                                            --
-- CERN BE-CO-HT         GN4124 core for PCIe FMC carrier                     --
--                       http://www.ohwr.org/projects/gn4124-core             --
--------------------------------------------------------------------------------
--
-- unit name: L2P_SER (l2p_ser.vhd)
--
-- author:
--
-- date:
--
-- version: 0.0
--
-- description: Generates the DDR L2P bus from SDR that is synchronous to ICLK
--
--
-- dependencies:
--
--------------------------------------------------------------------------------
-- last changes: <date> <initials> <log>
-- <extended description>
--------------------------------------------------------------------------------
-- TODO: -
--       -
--       -
--------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
use work.gn4124_core_pkg.all;


library UNISIM;
use UNISIM.vcomponents.all;

entity L2P_SER is
  port
    (
      ---------------------------------------------------------
      -- ICLK Clock Domain Inputs
      --
      ICLKp : in std_logic;
      ICLKn : in std_logic;
      IRST  : in std_logic;

      ICLK_VALID  : in  std_logic;
      ICLK_DFRAME : in  std_logic;
      ICLK_DATA   : in  std_logic_vector(31 downto 0);
      --
      ---------------------------------------------------------
      ---------------------------------------------------------
      -- SER Outputs
      --
      L2P_CLKp    : out std_logic;
      L2P_CLKn    : out std_logic;
      L2P_VALID   : out std_logic;
      L2P_DFRAME  : out std_logic;
      L2P_DATA    : out std_logic_vector(15 downto 0)
      --
      ---------------------------------------------------------
      );
end L2P_SER;

architecture BEHAVIOUR of L2P_SER is

-----------------------------------------------------------------------------
-- Internal Signals
-----------------------------------------------------------------------------
  signal ff_rst      : std_logic;
  signal Q_DFRAME    : std_logic;
  signal Q_VALID     : std_logic;
  signal Q_DATA      : std_logic_vector(ICLK_DATA'range);
  signal L2P_CLK_SDR : std_logic;


begin

  ------------------------------------------------------------------------------
  -- Active high reset for DDR FF
  ------------------------------------------------------------------------------
  gen_fifo_rst_n : if c_RST_ACTIVE = '0' generate
    ff_rst <= not(IRST);
  end generate;

  gen_fifo_rst : if c_RST_ACTIVE = '1' generate
    ff_rst <= IRST;
  end generate;


-----------------------------------------------------------------------------
-- Re-allign Data tightly for the +'ve clock edge
-----------------------------------------------------------------------------
  process (ICLKp, IRST)
  begin
    if(IRST = c_RST_ACTIVE) then
      Q_DFRAME <= '0';
      Q_VALID  <= '0';
      Q_DATA   <= (others => '0');
    elsif rising_edge(ICLKp) then
      Q_DFRAME <= ICLK_DFRAME;
      Q_VALID  <= ICLK_VALID;
      Q_DATA   <= ICLK_DATA;
    end if;
  end process;

  process (ICLKn, IRST)
  begin
    if(IRST = c_RST_ACTIVE) then
      L2P_VALID  <= '0';
      L2P_DFRAME <= '0';
    elsif rising_edge(ICLKn) then
      L2P_VALID  <= Q_VALID;
      L2P_DFRAME <= Q_DFRAME;
    end if;
  end process;


  DDROUT : for i in 0 to 15 generate
    U : OFDDRRSE
      port map
      (
        Q  => L2P_DATA(i),
        C0 => ICLKn,
        C1 => ICLKp,
        CE => '1',
        D0 => Q_DATA(i),
        D1 => Q_DATA(i+16),
        R  => ff_rst,
        S  => '0'
        );
  end generate;

  L2P_CLK_BUF : OBUFDS
    port map(
      O  => L2P_CLKp,
      OB => L2P_CLKn,
      I  => L2P_CLK_SDR);

  L2P_CLK_int : FDDRRSE
    port map(
      Q  => L2P_CLK_SDR,
      C0 => ICLKn,
      C1 => ICLKp,
      CE => '1',
      D0 => '1',
      D1 => '0',
      R  => '0',
      S  => '0');

end BEHAVIOUR;


