--------------------------------------------------------------------------------
--                                                                            --
-- CERN BE-CO-HT         GN4124 core for PCIe FMC carrier                     --
--                       http://www.ohwr.org/projects/gn4124-core             --
--------------------------------------------------------------------------------
--
-- unit name: 32 bit DMA master (l2p_dma_master.vhd)
--
-- author: Simon Deprez (simon.deprez@cern.ch)
--
-- date: 31-08-2010
--
-- version: 0.2
--
-- description: Provide a pipelined Wishbone interface to performs DMA
-- transfers from local application to PCI express host.
--
-- dependencies:
--
--------------------------------------------------------------------------------
-- last changes: <date> <initials> <log>
-- <extended description>
--------------------------------------------------------------------------------
-- TODO: - error signal
--       -
--       -
--------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;
use work.gn4124_core_pkg.all;


entity l2p_dma_master is
  port
    (
      ---------------------------------------------------------
      -- GN4124 core clock and reset
      sys_clk_i   : in std_logic;
      sys_rst_n_i : in std_logic;

      ---------------------------------------------------------
      -- From the DMA controller
      dma_ctrl_target_addr_i : in  std_logic_vector(31 downto 0);
      dma_ctrl_host_addr_h_i : in  std_logic_vector(31 downto 0);
      dma_ctrl_host_addr_l_i : in  std_logic_vector(31 downto 0);
      dma_ctrl_len_i         : in  std_logic_vector(31 downto 0);
      dma_ctrl_start_l2p_i   : in  std_logic;
      dma_ctrl_done_o        : out std_logic;
      dma_ctrl_error_o       : out std_logic;
      dma_ctrl_byte_swap_i   : in  std_logic_vector(1 downto 0);

      ---------------------------------------------------------
      -- To the L2P Interface (send the DMA data)
      ldm_arb_valid_o  : out std_logic;  -- Read completion signals
      ldm_arb_dframe_o : out std_logic;  -- Toward the arbiter
      ldm_arb_data_o   : out std_logic_vector(31 downto 0);
      ldm_arb_req_o    : out std_logic;
      arb_ldm_gnt_i    : in  std_logic;

      ---------------------------------------------------------
      -- DMA Interface (Pipelined Wishbone)
      l2p_dma_clk_i   : in  std_logic;                      -- Bus clock
      l2p_dma_adr_o   : out std_logic_vector(31 downto 0);  -- Adress
      l2p_dma_dat_i   : in  std_logic_vector(31 downto 0);  -- Data in
      l2p_dma_dat_o   : out std_logic_vector(31 downto 0);  -- Data out
      l2p_dma_sel_o   : out std_logic_vector(3 downto 0);   -- Byte select
      l2p_dma_cyc_o   : out std_logic;                      -- Read or write cycle
      l2p_dma_stb_o   : out std_logic;                      -- Read or write strobe
      l2p_dma_we_o    : out std_logic;                      -- Write
      l2p_dma_ack_i   : in  std_logic;                      -- Acknowledge
      l2p_dma_stall_i : in  std_logic                       -- for pipelined Wishbone
      );
end l2p_dma_master;


architecture behaviour of l2p_dma_master is

-----------------------------------------------------------------------------
-- Local constants
-----------------------------------------------------------------------------
  -- max payload set to 32 for debug/simul, should be 1024
  constant c_L2P_MAX_PAYLOAD      : unsigned(9 downto 0)         := to_unsigned(32, 10);
  signal   c_ADDR_FIFO_FULL_THRES : std_logic_vector(8 downto 0) := std_logic_vector(to_unsigned(500, 9));
  signal   c_DATA_FIFO_FULL_THRES : std_logic_vector(8 downto 0) := std_logic_vector(to_unsigned(500, 9));

-----------------------------------------------------------------------------
-- Internal Signals
-----------------------------------------------------------------------------
  -- Target address counter
  signal target_addr_cnt : unsigned(29 downto 0);
  signal dma_length_cnt  : unsigned(29 downto 0);

  -- Sync FIFOs
  signal fifo_rst        : std_logic;
  signal addr_fifo_rd    : std_logic;
  signal addr_fifo_valid : std_logic;
  signal addr_fifo_empty : std_logic;
  signal addr_fifo_dout  : std_logic_vector(31 downto 0);
  signal addr_fifo_din   : std_logic_vector(31 downto 0);
  signal addr_fifo_wr    : std_logic;
  signal addr_fifo_full  : std_logic;

  signal data_fifo_rd    : std_logic;
  signal data_fifo_valid : std_logic;
  signal data_fifo_empty : std_logic;
  signal data_fifo_dout  : std_logic_vector(31 downto 0);
  signal data_fifo_din   : std_logic_vector(31 downto 0);
  signal data_fifo_wr    : std_logic;
  signal data_fifo_full  : std_logic;

  -- Wishbone
  signal wb_read_cnt : unsigned(6 downto 0);
  signal wb_ack_cnt  : unsigned(6 downto 0);

  -- L2P DMA Master FSM
  type   l2p_dma_state_type is (IDLE, WB_DATA_WAIT, L2P_HEADER, L2P_ADDR_H, L2P_ADDR_L, L2P_DATA, L2P_DATA_LAST);
  signal l2p_dma_current_state : l2p_dma_state_type;

  -- L2P packet generator
  signal s_l2p_header : std_logic_vector(31 downto 0);
  signal s_l2p_data   : std_logic_vector(31 downto 0);

  signal l2p_len_cnt     : unsigned(29 downto 0);
  signal l2p_address_h   : unsigned(31 downto 0);
  signal l2p_address_l   : unsigned(31 downto 0);
  signal l2p_data_cnt    : unsigned(9 downto 0);
  signal l2p_64b_address : std_logic;

  signal l2p_byte_swap : std_logic_vector(1 downto 0);

begin


  ------------------------------------------------------------------------------
  -- Active high reset for fifo
  ------------------------------------------------------------------------------
  gen_fifo_rst_n : if c_RST_ACTIVE = '0' generate
    fifo_rst <= not(sys_rst_n_i);
  end generate;

  gen_fifo_rst : if c_RST_ACTIVE = '1' generate
    fifo_rst <= sys_rst_n_i;
  end generate;

  ------------------------------------------------------------------------------
  -- Target address counter
  ------------------------------------------------------------------------------
  p_target_cnt : process (sys_clk_i, sys_rst_n_i)
  begin
    if(sys_rst_n_i = c_RST_ACTIVE) then
      target_addr_cnt  <= (others => '0');
      dma_length_cnt   <= (others => '0');
      dma_ctrl_error_o <= '0';
      addr_fifo_wr     <= '0';
    elsif rising_edge(sys_clk_i) then
      if (dma_ctrl_start_l2p_i = '1') then
        if (l2p_dma_current_state = IDLE) then
          -- dma_ctrl_target_addr_i is a byte address and target_addr_cnt is a
          -- 32-bit word address
          target_addr_cnt  <= unsigned(dma_ctrl_target_addr_i(31 downto 2));
          -- dma_ctrl_len_i is in byte and dma_length_cnt is in 32-bit word
          dma_length_cnt   <= unsigned(dma_ctrl_len_i(31 downto 2));
          dma_ctrl_error_o <= '0';
        else
          target_addr_cnt  <= (others => '0');
          dma_length_cnt   <= (others => '0');
          dma_ctrl_error_o <= '1';
        end if;
      elsif (dma_length_cnt /= 0 and addr_fifo_full = '0') then
        addr_fifo_wr    <= '1';
        target_addr_cnt <= target_addr_cnt + 1;
        dma_length_cnt  <= dma_length_cnt - 1;
      else
        addr_fifo_wr <= '0';
      end if;
    end if;
  end process p_target_cnt;

  -- FIFO width is 32 bits
  addr_fifo_din <= "00" & std_logic_vector(target_addr_cnt);

  ------------------------------------------------------------------------------
  -- Packet generator
  ------------------------------------------------------------------------------
  -- Sends data to the host.
  -- Split in several packets if amont of data exceed max payload size.

  p_pkt_gen : process (sys_clk_i, sys_rst_n_i)
  begin
    if (sys_rst_n_i = c_RST_ACTIVE) then
      l2p_len_cnt     <= (others => '0');
      l2p_data_cnt    <= (others => '0');
      l2p_address_h   <= (others => '0');
      l2p_address_l   <= (others => '0');
      l2p_64b_address <= '0';
      l2p_byte_swap   <= (others => '0');
    elsif rising_edge(sys_clk_i) then
      -- First packet
      if (l2p_dma_current_state = IDLE) then
        if (dma_ctrl_start_l2p_i = '1') then
          l2p_len_cnt   <= unsigned(dma_ctrl_len_i(31 downto 2));
          l2p_address_h <= unsigned(dma_ctrl_host_addr_h_i);
          l2p_address_l <= unsigned(dma_ctrl_host_addr_l_i);
          l2p_byte_swap <= dma_ctrl_byte_swap_i;
        else
          if (l2p_len_cnt > c_L2P_MAX_PAYLOAD) then
            l2p_data_cnt <= c_L2P_MAX_PAYLOAD;
          else
            l2p_data_cnt <= l2p_len_cnt(9 downto 0);
          end if;
          if (l2p_address_h = 0) then
            l2p_64b_address <= '0';
          else
            l2p_64b_address <= '1';
          end if;
        end if;
        -- Next packet (if any)
      elsif (l2p_dma_current_state = L2P_ADDR_L) then
        if (l2p_len_cnt > c_L2P_MAX_PAYLOAD) then
          l2p_len_cnt <= l2p_len_cnt - c_L2P_MAX_PAYLOAD;
        else
          l2p_len_cnt <= (others => '0');
        end if;
      elsif (l2p_dma_current_state = L2P_DATA) then
        l2p_data_cnt <= l2p_data_cnt - 1;
      elsif (l2p_len_cnt > 0 and l2p_dma_current_state = L2P_DATA_LAST) then
        if (l2p_len_cnt > c_L2P_MAX_PAYLOAD) then
          l2p_data_cnt <= c_L2P_MAX_PAYLOAD;
        else
          l2p_data_cnt <= l2p_len_cnt(9 downto 0);
        end if;
      end if;
    end if;
  end process p_pkt_gen;

  -- Packet header
  s_l2p_header <= "000"                              -->  Traffic Class
                  & '0'                              -->  Snoop
                  & "001"                            -->  Memory write
                  & l2p_64b_address                  -->  Memory write
                  & "1111"                           -->  LBE
                  & "1111"                           -->  FBE
                  & "000"                            -->  Reserved
                  & '0'                              -->  VC
                  & "00"                             -->  Reserved
                  & std_logic_vector(l2p_data_cnt);  -->  Length

  -- Payload byte swap
  s_l2p_data <= data_fifo_dout when l2p_byte_swap = "00" else
                data_fifo_dout(15 downto 0)&
                data_fifo_dout(31 downto 16) when l2p_byte_swap = "10" else
                data_fifo_dout(7 downto 0)&
                data_fifo_dout(15 downto 8)&
                data_fifo_dout(23 downto 16)&
                data_fifo_dout(31 downto 24) when l2p_byte_swap = "11" else
                data_fifo_dout(23 downto 16)&
                data_fifo_dout(31 downto 24)&
                data_fifo_dout(7 downto 0)&
                data_fifo_dout(15 downto 8);

  -----------------------------------------------------------------------------
  -- L2P write FSM
  -----------------------------------------------------------------------------
  process(sys_clk_i, sys_rst_n_i)
  begin
    if (sys_rst_n_i = c_RST_ACTIVE) then
      l2p_dma_current_state <= IDLE;
      ldm_arb_req_o         <= '0';
      ldm_arb_data_o        <= (others => '0');
      ldm_arb_valid_o       <= '0';
      ldm_arb_dframe_o      <= '0';
      data_fifo_rd          <= '0';
      dma_ctrl_done_o       <= '0';
    elsif rising_edge(sys_clk_i) then
      case l2p_dma_current_state is
        -----------------------------------------------------------------
        -- IDLE
        -----------------------------------------------------------------
        when IDLE =>
          -- do nothing !
          data_fifo_rd     <= '0';
          dma_ctrl_done_o  <= '0';
          ldm_arb_data_o   <= (others => '0');
          ldm_arb_valid_o  <= '0';
          ldm_arb_dframe_o <= '0';

          if (data_fifo_empty = '0') then
            -- We have data to send -> prepare a packet, first the header
            l2p_dma_current_state <= L2P_HEADER;
            ldm_arb_req_o         <= '1';  -- request access to PCIe bus
            --ldm_arb_data_o        <= s_l2p_header;
            --ldm_arb_valid_o       <= '1';
            --ldm_arb_dframe_o      <= '1';
            --data_fifo_rd          <= '0';
            --dma_ctrl_done_o       <= '0';
            --else
            --l2p_dma_current_state <= IDLE;
          end if;

          -----------------------------------------------------------------
          -- L2P HEADER
          -----------------------------------------------------------------
        when L2P_HEADER =>
          if(arb_ldm_gnt_i = '1') then
            -- clear access request to the arbiter
            -- access is granted until dframe is cleared
            ldm_arb_req_o    <= '0';
            -- send header
            ldm_arb_data_o   <= s_l2p_header;
            ldm_arb_valid_o  <= '1';
            ldm_arb_dframe_o <= '1';
            if(l2p_64b_address = '1') then
              -- if host address is 64-bit, we have to send an additionnal
              -- 32-word containing highest bits of the host address
              l2p_dma_current_state <= L2P_ADDR_H;
              --ldm_arb_data_o        <= std_logic_vector(l2p_address_h);
              --ldm_arb_valid_o       <= '1';
              --ldm_arb_dframe_o      <= '1';
              --data_fifo_rd          <= '0';
            else
              -- for 32-bit host address, we only have to send lowest bits
              l2p_dma_current_state <= L2P_ADDR_L;
              -- Starts reading data in the fifo now, because there is
              -- 1 cycle delay until data are available
              data_fifo_rd          <= '1';
              --ldm_arb_data_o        <= std_logic_vector(l2p_address_l);
              --ldm_arb_valid_o       <= '1';
              --ldm_arb_dframe_o      <= '1';
            end if;
            --else
            --  l2p_dma_current_state <= L2P_HEADER;
            --  ldm_arb_req_o         <= '1';
            --  data_fifo_rd <= '0';
          end if;

          -----------------------------------------------------------------
          -- L2P ADDRESS (63-32)
          -----------------------------------------------------------------
        when L2P_ADDR_H =>
          -- send host address 32 highest bits
          ldm_arb_data_o        <= std_logic_vector(l2p_address_h);
          -- Now we still have to send lowest bits of the host address
          l2p_dma_current_state <= L2P_ADDR_L;
          -- Starts reading data in the fifo now, because there is
          -- 1 cycle delay until data are available
          data_fifo_rd          <= '1';
          --ldm_arb_data_o        <= std_logic_vector(l2p_address_l);
          --ldm_arb_valid_o       <= '1';
          --ldm_arb_dframe_o      <= '1';

          -----------------------------------------------------------------
          -- L2P ADDRESS (31-00)
          -----------------------------------------------------------------
        when L2P_ADDR_L =>
          -- send host address 32 lowest bits
          ldm_arb_data_o <= std_logic_vector(l2p_address_l);
          --if(data_fifo_valid = '1') then
          --  l2p_dma_current_state <= WB_DATA_WAIT;
          --  ldm_arb_valid_o       <= '0';
          --  ldm_arb_dframe_o      <= '1';
          --  data_fifo_rd          <= '1';
          if(l2p_data_cnt <= 2) then
            -- Only one 32-bit data word to send
            l2p_dma_current_state <= L2P_DATA_LAST;
            -- Stop reading from fifo
            data_fifo_rd          <= '0';
            --ldm_arb_data_o        <= s_l2p_data;
            --ldm_arb_valid_o       <= '1';
            --ldm_arb_dframe_o      <= '0';
          else
            -- More than one data word to send
            l2p_dma_current_state <= L2P_DATA;
            --ldm_arb_data_o <= s_l2p_data;
            --ldm_arb_valid_o       <= '0';
            --ldm_arb_dframe_o      <= '1';
            --if (data_fifo_empty = '0') then
            --  data_fifo_rd <= '1';
            --end if;
          end if;

          -----------------------------------------------------------------
          -- L2P DATA
          -----------------------------------------------------------------
        when L2P_DATA =>
          -- send data
          ldm_arb_data_o        <= s_l2p_data;
          ldm_arb_valid_o       <= '1';
          if(data_fifo_empty = '1') then
            l2p_dma_current_state <= WB_DATA_WAIT;
            --ldm_arb_valid_o       <= '0';
            --ldm_arb_dframe_o      <= '1';
            --data_fifo_rd          <= '1';
          elsif(l2p_data_cnt <= 2) then
            -- Only one 32-bit data word to send
            l2p_dma_current_state <= L2P_DATA_LAST;
            -- Stop reading from fifo
            data_fifo_rd          <= '0';
            --ldm_arb_data_o        <= s_l2p_data;
            --ldm_arb_valid_o       <= '1';
            --ldm_arb_dframe_o      <= '0';
          --else
          --  l2p_dma_current_state <= L2P_DATA;
          --  ldm_arb_data_o        <= s_l2p_data;
          --  ldm_arb_valid_o       <= '1';
          --  ldm_arb_dframe_o      <= '1';
          --  if (data_fifo_empty = '0') then
          --    data_fifo_rd <= '1';
          --  end if;
          end if;

          -----------------------------------------------------------------
          -- Wait data from the Wishbone machine
          -----------------------------------------------------------------
        when WB_DATA_WAIT =>
          ldm_arb_valid_o       <= '0';
          if(data_fifo_empty = '0') then
            l2p_dma_current_state <= L2P_DATA;
            --l2p_dma_current_state <= WB_DATA_WAIT;
            --ldm_arb_valid_o       <= '0';
            --ldm_arb_dframe_o      <= '1';
            --data_fifo_rd          <= '1';
          elsif(l2p_data_cnt <= 2) then
            -- Only one 32-bit data word to send
            l2p_dma_current_state <= L2P_DATA_LAST;
            -- Stop reading from fifo
            data_fifo_rd          <= '0';
            --ldm_arb_data_o        <= s_l2p_data;
            --ldm_arb_valid_o       <= '1';
            --ldm_arb_dframe_o      <= '0';
            --data_fifo_rd          <= '0';
          --else
          --  l2p_dma_current_state <= L2P_DATA;
          --  --ldm_arb_data_o <= s_l2p_data;
          --  ldm_arb_valid_o       <= '0';
          --  ldm_arb_dframe_o      <= '1';
          --  if (data_fifo_empty = '0') then
          --    data_fifo_rd <= '1';
          --  end if;
          end if;

          -----------------------------------------------------------------
          -- L2P DATA Last double word
          -----------------------------------------------------------------
        when L2P_DATA_LAST =>
          -- send the last data word
          ldm_arb_data_o        <= s_l2p_data;
          ldm_arb_valid_o       <= '1';
          -- clear dframe signal to indicate the end of packet
          ldm_arb_dframe_o      <= '0';
          if(l2p_len_cnt > 0) then
            -- There is still data to be send -> start a new packet
            l2p_dma_current_state <= L2P_HEADER;
            -- As the end of packet is used to delimit arbitration phases
            -- we have to ask again for permission
            ldm_arb_req_o         <= '1';
            --ldm_arb_data_o        <= s_l2p_header;
            --ldm_arb_valid_o       <= '1';
            --ldm_arb_dframe_o      <= '1';
            --data_fifo_rd          <= '0';
          else
            -- Nomore data to send, go back to sleep
            l2p_dma_current_state <= IDLE;
            -- Indicate that the DMA transfer is finished
            dma_ctrl_done_o       <= '1';
            --ldm_arb_data_o        <= (others => '0');
            --ldm_arb_valid_o       <= '0';
            --ldm_arb_dframe_o      <= '0';
            --data_fifo_rd          <= '0';
          end if;

          -----------------------------------------------------------------
          -- OTHERS
          -----------------------------------------------------------------
        when others =>
          -- should no arrive here, but just in case...
          l2p_dma_current_state <= IDLE;
          ldm_arb_req_o         <= '0';
          ldm_arb_data_o        <= (others => '0');
          ldm_arb_valid_o       <= '0';
          ldm_arb_dframe_o      <= '0';
          data_fifo_rd          <= '0';
          dma_ctrl_done_o       <= '0';

      end case;
    end if;
  end process;


--=========================================================================--
-- FIFOs for transition between GN4124 core and wishbone clock domain
--=========================================================================--
  cmp_addr_fifo : fifo_32x512
    port map (
      rst                     => fifo_rst,
      wr_clk                  => sys_clk_i,
      rd_clk                  => l2p_dma_clk_i,
      din                     => addr_fifo_din,
      wr_en                   => addr_fifo_wr,
      rd_en                   => addr_fifo_rd,
      prog_full_thresh_assert => c_ADDR_FIFO_FULL_THRES,
      prog_full_thresh_negate => c_ADDR_FIFO_FULL_THRES,
      dout                    => addr_fifo_dout,
      full                    => open,
      empty                   => addr_fifo_empty,
      valid                   => addr_fifo_valid,
      prog_full               => addr_fifo_full);

  cmp_data_fifo : fifo_32x512
    port map (
      rst                     => fifo_rst,
      wr_clk                  => l2p_dma_clk_i,
      rd_clk                  => sys_clk_i,
      din                     => data_fifo_din,
      wr_en                   => data_fifo_wr,
      rd_en                   => data_fifo_rd,
      prog_full_thresh_assert => c_DATA_FIFO_FULL_THRES,
      prog_full_thresh_negate => c_DATA_FIFO_FULL_THRES,
      dout                    => data_fifo_dout,
      full                    => open,
      empty                   => data_fifo_empty,
      valid                   => data_fifo_valid,
      prog_full               => data_fifo_full);

  data_fifo_din <= l2p_dma_dat_i;
  data_fifo_wr  <= l2p_dma_ack_i;

--=========================================================================--
-- Pipelined wishbone master
--=========================================================================--
-- Initatiates read transactions as long there is an address present
-- in the address fifo. Then fills the data fifo with the read data.

  -- Wishbone master only make reads
  l2p_dma_we_o  <= '0';
  l2p_dma_dat_o <= (others => '0');

  -- Read address FIFO
  addr_fifo_rd <= not(addr_fifo_empty)
                  and not(l2p_dma_stall_i)
                  and not(data_fifo_full);

  -- Wishbone master process
  p_wb_master : process (l2p_dma_clk_i, sys_rst_n_i)
  begin
    if (sys_rst_n_i = c_RST_ACTIVE) then
      l2p_dma_adr_o <= (others => '0');
      l2p_dma_stb_o <= '0';
      l2p_dma_cyc_o <= '0';
      l2p_dma_sel_o <= (others => '0');
    elsif rising_edge(l2p_dma_clk_i) then
      -- adr
      if (addr_fifo_valid = '1') then
        l2p_dma_adr_o <= addr_fifo_dout;
      end if;
      -- stb and sel
      if (addr_fifo_valid = '1' or l2p_dma_stall_i = '1') then
        l2p_dma_stb_o <= '1';
        l2p_dma_sel_o <= (others => '1');
      else
        l2p_dma_stb_o <= '0';
        l2p_dma_sel_o <= (others => '0');
      end if;
      -- cyc
      if (addr_fifo_valid = '1') then
        l2p_dma_cyc_o <= '1';
      elsif (wb_ack_cnt-1 = wb_read_cnt and l2p_dma_ack_i = '1') then
        l2p_dma_cyc_o <= '0';
      end if;
    end if;
  end process p_wb_master;

  -- Wishbone read cycle counter
  p_wb_read_cnt : process (l2p_dma_clk_i, sys_rst_n_i)
  begin
    if (sys_rst_n_i = c_RST_ACTIVE) then
      wb_read_cnt <= (others => '0');
    elsif rising_edge(l2p_dma_clk_i) then
      if (addr_fifo_valid = '1') then
        wb_read_cnt <= wb_read_cnt + 1;
      end if;
    end if;
  end process p_wb_read_cnt;

-- Wishbone ack counter
  p_wb_ack_cnt : process (l2p_dma_clk_i, sys_rst_n_i)
  begin
    if (sys_rst_n_i = c_RST_ACTIVE) then
      wb_ack_cnt <= (others => '0');
    elsif rising_edge(l2p_dma_clk_i) then
      if (l2p_dma_ack_i = '1') then
        wb_ack_cnt <= wb_ack_cnt + 1;
      end if;
    end if;
  end process p_wb_ack_cnt;


end behaviour;

